LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY conv_7seg IS
PORT (D:IN STD_LOGIC_VECTOR(3 DOWNTO 0);
O:OUT STD_LOGIC_VECTOR(6 DOWNTO 0));
END conv_7seg;
ARCHITECTURE RTL OF conv_7seg IS
BEGIN
PROCESS (D)
BEGIN
CASE D IS
WHEN "0000"=>O<="1111110";
WHEN "0001"=>O<="0110000";
WHEN "0010"=>O<="1101101";
WHEN "0011"=>O<="1111001";
WHEN "0100"=>O<="0110011";
WHEN "0101"=>O<="1011011";
WHEN "0110"=>O<="0011111";
WHEN "0111"=>O<="1110000";
WHEN "1000"=>O<="1111111";
WHEN "1001"=>O<="1110011";
WHEN OTHERS=>O<="XXXXXXX";
END CASE;
END PROCESS;
END RTL;