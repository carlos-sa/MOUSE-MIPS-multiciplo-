LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY conv_7seg IS
PORT (D:IN STD_LOGIC_VECTOR(3 DOWNTO 0);
O:OUT STD_LOGIC_VECTOR(6 DOWNTO 0));
END conv_7seg;
ARCHITECTURE RTL OF conv_7seg IS
BEGIN
PROCESS (D)
BEGIN
CASE D IS
WHEN "0000"=>O<="0000001";
WHEN "0001"=>O<="1001111";
WHEN "0010"=>O<="0010010";
WHEN "0011"=>O<="0000110";
WHEN "0100"=>O<="1001100";
WHEN "0101"=>O<="0100100";
WHEN "0110"=>O<="1100000";
WHEN "0111"=>O<="0001111";
WHEN "1000"=>O<="0000000";
WHEN "1001"=>O<="0001100";
WHEN OTHERS=>O<="XXXXXXX";
END CASE;
END PROCESS;
END RTL;